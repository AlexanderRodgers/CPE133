`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 05/10/2019 11:06:00 AM
// Design Name: 
// Module Name: 4bit_Dcom
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module 4bit_Dcom(
    input [3:0] D,
    input clk,
    input clr,
    input set,
    output [3:0] Q
    );
endmodule
