module JKFF(input clr, input clk, input [1:0] JK, output reg Q, output Qb);
assign Qb=~Q;
always @(posedge clk)
  if (clr) Q<=1'b0; else
  case (JK)
 2'b00: Q<=Q;
 2'b01: Q<=1'b0;
 2'b10: Q<=1'b1;
 2'b11: Q<=~Q;
 endcase
endmodule